library verilog;
use verilog.vl_types.all;
entity electronic_enigma_vlg_vec_tst is
end electronic_enigma_vlg_vec_tst;
